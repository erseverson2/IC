module pielineIF(clk,rst,,,);


Register_4_Bit( input clk, input rst, input [3:0] D, input WriteReg, input ReadEnable1, input ReadEnable2, inout [3:0] Bitline1, inout [3:0] Bitline2);
Register_4_Bit( input clk, input rst, input [3:0] D, input WriteReg, input ReadEnable1, input ReadEnable2, inout [3:0] Bitline1, inout [3:0] Bitline2);
Register_4_Bit( input clk, input rst, input [3:0] D, input WriteReg, input ReadEnable1, input ReadEnable2, inout [3:0] Bitline1, inout [3:0] Bitline2);


endmodule