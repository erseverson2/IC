module pielineMEM(,,,,);



dff (q, d, wen, clk, rst);
Register(input clk, input rst, input [15:0] D, input WriteReg, input ReadEnable1, input ReadEnable2, inout [15:0] Bitline1, inout [15:0] Bitline2);



endmodule